---------------------------------------------------------------------------
-- control_unit.vhd - Control Unit Implementation
--
-- Notes: refer to headers in single_cycle_core.vhd for the supported ISA.
--
--  control signals:
--     reg_dst    : asserted for ADD instructions, so that the register
--                  destination number for the 'write_register' comes from
--                  the rd field (bits 3-0). 
--     reg_write  : asserted for ADD and LOAD instructions, so that the
--                  register on the 'write_register' input is written with
--                  the value on the 'write_data' port.
--     alu_src    : asserted for LOAD and STORE instructions, so that the
--                  second ALU operand is the sign-extended, lower 4 bits
--                  of the instruction.
--     mem_write  : asserted for STORE instructions, so that the data 
--                  memory contents designated by the address input are
--                  replaced by the value on the 'write_data' input.
--     mem_to_reg : asserted for LOAD instructions, so that the value fed
--                  to the register 'write_data' input comes from the
--                  data memory.
--
--
-- Copyright (C) 2006 by Lih Wen Koh (lwkoh@cse.unsw.edu.au)
-- All Rights Reserved. 
--
-- The single-cycle processor core is provided AS IS, with no warranty of 
-- any kind, express or implied. The user of the program accepts full 
-- responsibility for the application of the program and the use of any 
-- results. This work may be downloaded, compiled, executed, copied, and 
-- modified solely for nonprofit, educational, noncommercial research, and 
-- noncommercial scholarship purposes provided that this notice in its 
-- entirety accompanies all copies. Copies of the modified software can be 
-- delivered to persons who use it solely for nonprofit, educational, 
-- noncommercial research, and noncommercial scholarship purposes provided 
-- that this notice in its entirety accompanies all copies.
--
---------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity control_unit is
    port ( opcode     : in  std_logic_vector(3 downto 0);
           --reg_dst    : out std_logic;
           reg_write  : out std_logic;
           alu_src    : out std_logic;
			  beq			 : out std_logic;
           mem_write  : out std_logic;
           alu_ctrl   : out std_logic_vector(3 downto 0);
           mem_to_reg : out std_logic; 
			  jmp        : out std_logic);
end control_unit;

architecture behavioural of control_unit is
			
constant OP_AND   : std_logic_vector(3 downto 0) := "0000";
constant OP_ANDI  : std_logic_vector(3 downto 0) := "0001";
constant OP_XOR   : std_logic_vector(3 downto 0) := "0010";
constant OP_ADD   : std_logic_vector(3 downto 0) := "0011";
constant OP_ADDI  : std_logic_vector(3 downto 0) := "0100";
constant OP_LW    : std_logic_vector(3 downto 0) := "0101";
constant OP_SWI   : std_logic_vector(3 downto 0) := "0110";
constant OP_SRLI  : std_logic_vector(3 downto 0) := "0111";
constant OP_SRL   : std_logic_vector(3 downto 0) := "1000";
constant OP_SLLI  : std_logic_vector(3 downto 0) := "1001";
constant OP_BEQ   : std_logic_vector(3 downto 0) := "1010";
constant OP_JUMP  : std_logic_vector(3 downto 0) := "1011";
--constant OP_SLT   : std_logic_vector(3 downto 0) := "1100";
constant OP_J     : std_logic_vector(3 downto 0) := "1110";

begin

	--high when its a sub
    alu_ctrl(3)   <= '1' when (opcode = OP_BEQ) else
							'0';
							
	 alu_ctrl(2)	<= '0' when (opcode = OP_SLLI) else
							'1';
							
	 alu_ctrl(1)	<= '0' when (opcode = OP_AND
										 or opcode = OP_ANDI
										 or opcode = OP_XOR) else
							'1';
							
	 alu_ctrl(0)	<= '1' when (opcode = OP_AND
										 or opcode = OP_ANDI
										 or opcode = OP_SRLI
										 or opcode = OP_SRL
										 or opcode = OP_SLLI) else
							'0';

    --reg_dst    <= '1' when opcode = OP_ADD else
    --              '0';

	 jmp			<= '1' when (opcode = OP_JUMP) else
						'0';

	 beq			<= '1' when (opcode = OP_BEQ) else
						'0';

    reg_write  <= '0' when (opcode = OP_SWI 
                            or opcode = OP_BEQ
									 or opcode = OP_JUMP) else
                  '1';
    
	 --for usage of immediates
    alu_src    <= '1' when (opcode = OP_ANDI 
                           or opcode = OP_ADDI
									or opcode = OP_SWI
									--or opcode = OP_LW
									or opcode = OP_SRLI
									or opcode = OP_SLLI) else
                  '0';
                 
    mem_write  <= '1' when (opcode = OP_SWI) else
                  '0';
                 
    mem_to_reg <= '1' when opcode = OP_LW else
                  '0';

end behavioural;
